library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;

library std;
use std.textio.all;

entity data_maker is
  port (
    CLK  : in  std_logic;
    RST_n   : in  std_logic;
    VOUT    : out std_logic;
    DOUT : out std_logic_vector(31 downto 0);
    END_SIM : out std_logic);
end data_maker;

architecture beh of data_maker is

  constant tco : time := 1 ns;

  signal sEndSim: std_logic;
  signal END_SIM_i: std_logic_vector(0 to 5);

begin  -- beh

  process (CLK, RST_n)
    file fp : text open read_mode is "C:\Users\nicola\OneDrive\Desktop\ISA\ISAL2\tb\fp_samples.hex";
    variable ptr : line;
    variable val : std_logic_vector(31 downto 0);
  begin  -- process
    if RST_n = '0' then                 -- asynchronous reset (active low)
      DOUT <= (others => '0') after tco;      
      VOUT <= '0' after tco;
      sEndSim <= '0' after tco;
    elsif CLK'event and CLK = '1' then  -- rising clock edge
      if (not(endfile(fp))) then
        readline(fp, ptr);
        hread(ptr, val);
        DOUT <= val after tco;
        VOUT <= '1' after tco;
        sEndSim <= '0' after 5*tco;
      else
        VOUT <= '0' after tco;        
        sEndSim <= '1' after tco;
      end if;
    end if;
  end process;

  process (CLK, RST_n)
  begin  -- process
    if RST_n = '0' then                 -- asynchronous reset (active low)
      END_SIM_i <= (others => '0') after tco;
    elsif CLK'event and CLK = '1' then  -- rising clock edge
      END_SIM_i(0) <= sEndSim after tco;
      END_SIM_i   (1 to 5) <= END_SIM_i(0 to 4) after tco;
    end if;
  end process;

  END_SIM <= END_SIM_i(5); 

end beh;
